// Request-Grant-Done arbiter as describe pages 213/215 of 
// Synchronization and Arbitration in Digital Systems
//   Author:	David J. Kinniment
// Wiley Publishing ©2008 
// ISBN:047051082X 9780470510827


module rgd_arbitrer(/*AUTOARG*/
   // Outputs
   g1, g2,
   // Inputs
   r1, d1, r2, d2, rstn
   );
   input r1;
   input d1;
   input r2;
   input d2;
   output g1;
   output g2;

   input  rstn;
   
   



endmodule // rgd_arbitrer

